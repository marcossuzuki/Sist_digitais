library verilog;
use verilog.vl_types.all;
entity somador_paralelo_4bits_vlg_vec_tst is
end somador_paralelo_4bits_vlg_vec_tst;
