library verilog;
use verilog.vl_types.all;
entity bcd_behavioral_vlg_check_tst is
    port(
        Bv              : in     vl_logic_vector(7 downto 0);
        sampler_rx      : in     vl_logic
    );
end bcd_behavioral_vlg_check_tst;
