library verilog;
use verilog.vl_types.all;
entity somador_completo_vlg_vec_tst is
end somador_completo_vlg_vec_tst;
