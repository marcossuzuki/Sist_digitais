library verilog;
use verilog.vl_types.all;
entity somador_bin_par_vlg_vec_tst is
end somador_bin_par_vlg_vec_tst;
