library verilog;
use verilog.vl_types.all;
entity mux_4_1_vlg_check_tst is
    port(
        F0              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux_4_1_vlg_check_tst;
