library verilog;
use verilog.vl_types.all;
entity decoder_BCD_7seg_vlg_vec_tst is
end decoder_BCD_7seg_vlg_vec_tst;
