library verilog;
use verilog.vl_types.all;
entity mux_2_1_vlg_check_tst is
    port(
        F               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux_2_1_vlg_check_tst;
